library ieee;
use ieee.std_logic_1164.all;

entity bloqueio_ula is
	port(
        s_block : in std_logic;
        s_in    : in std_logic;

        s    : out std_logic  
	);
end bloqueio_ula;

architecture comp of porta_AND_8in is
    begin
        


end architecture;