library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity ULA is
	port(
        cac      : in std_logic_vector(7 downto 0);

	);
end ULA;
